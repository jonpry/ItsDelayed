.title KiCad schematic



.func E(x) {exp(x)}

.include "ff_nonfet.cor"

*.include "lod_params.cor"

***************************************************
*                RO DLC FACTORS                   *
***************************************************
.param
+ lv_dlc_rotweak               = 00.00e-9
+ lvhvt_dlc_rotweak            = 00.00e-9
+ lvt_dlc_rotweak              = 00.00e-9
+ hv_dlc_rotweak               =  00.00e-9
+ nshort_dlc_rotweak           =  lv_dlc_rotweak
+ nshortesd_dlc_rotweak        =  lv_dlc_rotweak
+ nlowvt_dlc_rotweak           =  lvt_dlc_rotweak
+ pshort_dlc_rotweak           =  lv_dlc_rotweak
+ plowvt_dlc_rotweak           =  lvt_dlc_rotweak
+ phighvt_dlc_rotweak          =  lvhvt_dlc_rotweak
+ nhvesd_dlc_rotweak           =  hv_dlc_rotweak
+ phvesd_dlc_rotweak           =  hv_dlc_rotweak
+ ntvnative_dlc_rotweak        =  hv_dlc_rotweak
+ nhvnative_dlc_rotweak        =  hv_dlc_rotweak
+ nhv_dlc_rotweak              =  hv_dlc_rotweak
+ phv_dlc_rotweak              =  hv_dlc_rotweak
+ pvhv_dlc_rotweak              =  hv_dlc_rotweak
*
+ npass_dlc_rotweak            =  lv_dlc_rotweak
+ npassll_dlc_rotweak          =  lv_dlc_rotweak
+ fnpass_dlc_rotweak           =  hv_dlc_rotweak
+ npd_dlc_rotweak              =  lv_dlc_rotweak
+ npdll_dlc_rotweak            =  lv_dlc_rotweak
+ ppu_dlc_rotweak              =  lv_dlc_rotweak
+ ppull_dlc_rotweak            =  lv_dlc_rotweak
*
+ sonos_e_dlc_rotweak          =  hv_dlc_rotweak
+ sonos_p_dlc_rotweak          =  hv_dlc_rotweak
+ sonos_eeol_dlc_rotweak       =  hv_dlc_rotweak
+ sonos_peol_dlc_rotweak       =  hv_dlc_rotweak


.include nlowvt_mm.cor
.include nlowvt_ff.cor
.include nlowvt.pm3

.include pshort_mm.cor
.include pshort_ff.cor
.include pshort.pm3

.option scale=1U
.include TOP.spice

*.subckt TOP S SB VSS VDD OUT0 OUT OUT2 OUT3 OUT4 OUT5 OUT6 S4B S4 S2B S2 S3B S3 OUTD IN OUT OUTDD OUTDDD
*.subckt TOP S SB VSS VDD OUT0 OUT OUT2 OUT3 OUT4 OUT5 OUT6 S4B S4 S2B S2 S3B S3 OUTD IN OUT OUTDD OUTDDD
*.subckt TOP S SB VSS VDD S4B S4 S2B S2 S3B S3 OUTD IN OUT OUTDD OUTDDD
*.subckt TOP S SB VSS VDD OUT7 S2B S2 S3B S3 S4B S4 OUTD IN OUT OUTDD OUTDDD OUTDDDD
*.subckt TOP S SB VSS VDD S2B S2 S3B S3 S4B S4 S5B S5 OUTD IN OUT OUTDD OUTDDD OUTDDDD
*.subckt TOP S SB VSS VDD S2B S2 S3B S3 S4B S4 S5B S5 OUTD IN OUT OUTDDDDD OUTDD OUTDDD OUTDDDD
*.SUBCKT TOP VSS IN OUTDDDDD OUTD OUT OUTDD OUTDDD OUTDDDD S5 S5B SB S VDD S2 S2B S3 S3B S4 S4B

   
X1 gnd IN OUTDDDDD OUTD OUT OUTDD OUTDDD OUTDDDD ctrl5 ctrl5b ctrlb ctrl pwr ctrl2 ctrl2b ctrl3 ctrl3b ctrl4 ctrl4b TOP
Vpos pwr gnd DC 1.8V 
Vctrl ctrl gnd DC 1.8V 
Vctrlb ctrlb gnd DC 0V 
Vctrl2 ctrl2 gnd DC 1.8V 
Vctrl2b ctrl2b gnd DC 0V
Vctrl3 ctrl3 gnd DC 0V       
Vctrl3b ctrl3b gnd DC 1.8V  
Vctrl4 ctrl4 gnd DC 0V       
Vctrl4b ctrl4b gnd DC 1.8V  
Vctrl5 ctrl5 gnd DC 1.8V       
Vctrl5b ctrl5b gnd DC 0V  
Vsig in2 gnd DC 0V PULSE(0 1.8V 0 100p 100p 500p 1n) 
R10001 in in2 1k


*.OPTION ABSTOL=1e-15.
*.OPTION GMIN=1.0e-10.
*.OPTION ITL1=1e5
*.OPTION RSHUNT=1e12
*.OPTION RELTOL=1e-5
*.op
.control
TRAN 10p 5N
alter @Vctrl[dc] = 0V
alter @Vctrlb[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl2[dc] = 0V
alter @Vctrl2b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl[dc] = 1.8V
alter @Vctrlb[dc] = 0V
TRAN 10p 5N
alter @Vctrl2[dc] = 1.8V
alter @Vctrl2b[dc] = 0V
TRAN 10p 5N
alter @Vctrl3[dc] = 1.8V
alter @Vctrl3b[dc] = 0V
TRAN 10p 5N
alter @Vctrl[dc] = 0V
alter @Vctrlb[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl2[dc] = 0V
alter @Vctrl2b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl[dc] = 1.8V
alter @Vctrlb[dc] = 0V
TRAN 10p 5N
alter @Vctrl2[dc] = 1.8V
alter @Vctrl2b[dc] = 0V
TRAN 10p 5N
alter @Vctrl3[dc] = 0V
alter @Vctrl3b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl4[dc] = 1.8V
alter @Vctrl4b[dc] = 0V
TRAN 10p 5N
alter @Vctrl[dc] = 0V
alter @Vctrlb[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl2[dc] = 0V
alter @Vctrl2b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl[dc] = 1.8V
alter @Vctrlb[dc] = 0V
TRAN 10p 5N
alter @Vctrl2[dc] = 1.8V
alter @Vctrl2b[dc] = 0V
TRAN 10p 5N
alter @Vctrl3[dc] = 1.8V
alter @Vctrl3b[dc] = 0V
TRAN 10p 5N
alter @Vctrl[dc] = 0V
alter @Vctrlb[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl2[dc] = 0V
alter @Vctrl2b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl[dc] = 1.8V
alter @Vctrlb[dc] = 0V
TRAN 10p 5N
alter @Vctrl2[dc] = 1.8V
alter @Vctrl2b[dc] = 0V
TRAN 10p 5N
alter @Vctrl3[dc] = 0V
alter @Vctrl3b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl5[dc] = 0V
alter @Vctrl5b[dc] = 1.8V
alter @Vctrl4[dc] = 0V
alter @Vctrl4b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl[dc] = 0V
alter @Vctrlb[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl2[dc] = 0V
alter @Vctrl2b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl[dc] = 1.8V
alter @Vctrlb[dc] = 0V
TRAN 10p 5N
alter @Vctrl2[dc] = 1.8V
alter @Vctrl2b[dc] = 0V
TRAN 10p 5N
alter @Vctrl3[dc] = 1.8V
alter @Vctrl3b[dc] = 0V
TRAN 10p 5N
alter @Vctrl[dc] = 0V
alter @Vctrlb[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl2[dc] = 0V
alter @Vctrl2b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl[dc] = 1.8V
alter @Vctrlb[dc] = 0V
TRAN 10p 5N
alter @Vctrl2[dc] = 1.8V
alter @Vctrl2b[dc] = 0V
TRAN 10p 5N
alter @Vctrl3[dc] = 0V
alter @Vctrl3b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl4[dc] = 1.8V
alter @Vctrl4b[dc] = 0V
TRAN 10p 5N
alter @Vctrl[dc] = 0V
alter @Vctrlb[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl2[dc] = 0V
alter @Vctrl2b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl[dc] = 1.8V
alter @Vctrlb[dc] = 0V
TRAN 10p 5N
alter @Vctrl2[dc] = 1.8V
alter @Vctrl2b[dc] = 0V
TRAN 10p 5N
alter @Vctrl3[dc] = 1.8V
alter @Vctrl3b[dc] = 0V
TRAN 10p 5N
alter @Vctrl[dc] = 0V
alter @Vctrlb[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl2[dc] = 0V
alter @Vctrl2b[dc] = 1.8V
TRAN 10p 5N
alter @Vctrl[dc] = 1.8V
alter @Vctrlb[dc] = 0V
TRAN 10p 5N
alter @Vctrl2[dc] = 1.8V
alter @Vctrl2b[dc] = 0V
TRAN 10p 5N
alter @Vctrl3[dc] = 0V
alter @Vctrl3b[dc] = 1.8V
TRAN 10p 5N

plot v(in) tran2.v(outddddd) tran3.v(outddddd) tran4.v(outddddd) tran5.v(outddddd) tran6.v(outddddd) tran7.v(outddddd) tran8.v(outddddd) tran9.v(outddddd) tran10.v(outddddd) tran11.v(outddddd) tran12.v(outddddd) tran13.v(outddddd) tran14.v(outddddd) tran15.v(outddddd) tran16.v(outddddd) tran17.v(outddddd) tran18.v(outddddd) tran19.v(outddddd) tran20.v(outddddd) tran21.v(outddddd) tran22.v(outddddd) tran23.v(outddddd) tran24.v(outddddd) tran25.v(outddddd) tran26.v(outddddd) tran27.v(outddddd) tran28.v(outddddd) tran29.v(outddddd) tran30.v(outddddd) tran31.v(outddddd) tran32.v(outddddd) tran33.v(outddddd) tran34.v(outddddd) tran35.v(outddddd) tran36.v(outddddd) tran37.v(outddddd) tran38.v(outddddd) tran39.v(outddddd) tran40.v(outddddd) tran41.v(outddddd) tran42.v(outddddd) tran43.v(outddddd)

*plot v(in) tran6.v(outddd) tran7.v(outddd) tran8.v(outddd) tran9.v(outddd)
*plot v(in) v(out0) v(out) v(out2) v(out3) v(out4) v(out5) v(out6)

*plot v(in) v(outddd)

.endc

.end
